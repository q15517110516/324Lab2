library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity Mux_tb is
--  Port ( );
end Mux_tb;

architecture Behavioral of Mux_tb is
component mux4
    port( 
      i0 : in std_logic;
      i1 : in std_logic;
      i2 : in std_logic;
      i3 : in std_logic;
      sel: in std_logic_vector(1 downto 0);
      o  : out std_logic);
end component;
signal i0,i1,i2,i3,o : std_logic;
signal sel:std_logic_vector(1 downto 0);
begin
mux4_0: mux4 port map (i0=>i0,i1=>i1,i2=>i2,i3=>i3,sel=>sel,o=>o);
process
type pat_type is record
i0,i1,i2,i3:std_logic;
sel:std_logic_vector(1 downto 0);
o:std_logic;
end record;
type pat_arr is array (natural range<>) of pat_type;
constant pat : pat_arr:=
(
    ('0','0','0','0',"00",'0'),			--data format is  i0  i1   i2   i3   sel   o
    ('0','0','0','0',"01",'0'),
    ('0','0','0','0',"11",'0'),
    ('0','0','0','0',"10",'0'),
    
    ('0','0','0','1',"00",'1'),
    ('0','0','0','1',"01",'0'),
    ('0','0','0','1',"11",'0'),
    ('0','0','0','1',"10",'0'),
    
    ('0','0','1','0',"00",'0'),
    ('0','0','1','0',"01",'1'),
    ('0','0','1','0',"11",'0'),
    ('0','0','1','0',"10",'0'),
    
    ('0','0','1','1',"00",'1'),
    ('0','0','1','1',"01",'1'),
    ('0','0','1','1',"11",'0'),
    ('0','0','1','1',"10",'0'),
    
    ('0','1','0','0',"00",'0'),
    ('0','1','0','0',"01",'0'),
    ('0','1','0','0',"11",'1'),
    ('0','1','0','0',"10",'0'),

    ('0','1','0','1',"00",'1'),
    ('0','1','0','1',"01",'0'),
    ('0','1','0','1',"11",'1'),
    ('0','1','0','1',"10",'0'),

    ('0','1','1','0',"00",'0'),
    ('0','1','1','0',"01",'1'),
    ('0','1','1','0',"11",'1'),
    ('0','1','1','0',"10",'0'),
    
    ('0','1','1','1',"00",'1'),
    ('0','1','1','1',"01",'1'),
    ('0','1','1','1',"11",'1'),
    ('0','1','1','1',"10",'0'),

    ('1','0','0','0',"00",'0'),
    ('1','0','0','0',"01",'0'),
    ('1','0','0','0',"11",'0'),
    ('1','0','0','0',"10",'1'),
  
    ('1','0','0','1',"00",'1'),
    ('1','0','0','1',"01",'0'),
    ('1','0','0','1',"11",'0'),
    ('1','0','0','1',"10",'1'),

    ('1','0','0','1',"00",'1'),
    ('1','0','0','1',"01",'0'),
    ('1','0','0','1',"11",'0'),
    ('1','0','0','1',"10",'1'),

    ('1','0','1','0',"00",'0'),
    ('1','0','1','0',"01",'1'),
    ('1','0','1','0',"11",'0'),
    ('1','0','1','0',"10",'1'),
    
    ('1','0','1','1',"00",'1'),
    ('1','0','1','1',"01",'1'),
    ('1','0','1','1',"11",'0'),
    ('1','0','1','1',"10",'1'),

    ('1','1','0','0',"00",'0'),
    ('1','1','0','0',"01",'0'),
    ('1','1','0','0',"11",'1'),
    ('1','1','0','0',"10",'1'),

    ('1','1','0','1',"00",'1'),
    ('1','1','0','1',"01",'0'),
    ('1','1','0','1',"11",'1'),
    ('1','1','0','1',"10",'1'),
    
    ('1','1','1','0',"00",'0'),
    ('1','1','1','0',"01",'1'),
    ('1','1','1','0',"11",'1'),
    ('1','1','1','0',"10",'1'),
    
    ('1','1','1','1',"00",'1'),
    ('1','1','1','1',"01",'1'),
    ('1','1','1','1',"11",'1'),
    ('1','1','1','1',"10",'1')
);
begin
    for n in pat'range loop
    i0<=pat(n).i0;
    i1<=pat(n).i1;
    i2<=pat(n).i2;
    i3<=pat(n).i3;
    sel<=pat(n).sel;
    wait for 10ns;
    
    assert o<=pat(n).o 
    report "bad output value" severity error;
 end loop;
assert false report "end of test" severity note;
wait;

end process;
end Behavioral;
